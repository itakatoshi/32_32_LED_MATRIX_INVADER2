
module opening (
    input clk,
    input reset,
    input wire [4:0] col,
    input wire [3:0] row,
    input wire sw0_raise,
    input wire sw1_raise,
    input wire sw2_raise,
    input wire sw3_raise,
    input wire [2:0]cur_stage,
    output reg sound_en,
    //output reg [3:0] note_sel,
    output wire [2:0]next_stage_flag,
    output wire [1:0] stage_select,
    output wire RED_UP_WIRE,
    output wire RED_DOWN_WIRE,
    output wire GREEN_UP_WIRE,
    output wire GREEN_DOWN_WIRE
//    output wire BLUE_UP_WIRE,
//    output wire BLUE_DOWN_WIRE
);

// ��Ԃ������萔���`
parameter OPENING = 3'b000;
parameter STAGE1  = 3'b001;
parameter STAGE2  = 3'b010;
parameter STAGE3  = 3'b011;
parameter FINISH  = 3'b100;

//���d�u�U�[�̐���
reg [2:0] next_stage;
reg [1:0] stage_select_flag; 

// 2������ reg �z��
reg [31:0] R_UP [15:0], R_DOWN [15:0], G_UP [15:0], G_DOWN [15:0]; //B_UP [15:0], B_DOWN [15:0];
reg [23:0] count;
reg [23:0] MAX;

// �u�U�[�J�E���g
reg [16:0]sound_count;
parameter BOM_SOUND = 81_250; //12MHz  


assign RED_UP_WIRE = R_UP[row][col];
assign RED_DOWN_WIRE = R_DOWN[row][col];
assign GREEN_UP_WIRE = G_UP[row][col];
assign GREEN_DOWN_WIRE = G_DOWN[row][col];
//assign BLUE_UP_WIRE = B_UP[row][col];
//assign BLUE_DOWN_WIRE = B_DOWN[row][col];
assign stage_select = stage_select_flag;
assign next_stage_flag = next_stage;



always @(posedge clk or posedge reset) begin
    
    
	if(reset) begin
	
        G_UP[0]<=32'b11111111111111111111111111111111;
        G_UP[1]<=32'b10000000000000000000000000000001;
        G_UP[2]<=32'b10000000000000000000000000000001;
        G_UP[3]<=32'b10000000000000000000000000000001;
        G_UP[4]<=32'b10000000000000000000000000000001;
        G_UP[5]<=32'b10111111110001000010000001100001;
        G_UP[6]<=32'b10111111110000100100000011110001;
        G_UP[7]<=32'b10111111110010111101000111111001;
        G_UP[8]<=32'b10111111110011011011001101101101;
        G_UP[9]<=32'b10111111110011111111001111111101;
        G_UP[10]<=32'b10111111110001111110000010010001;
        G_UP[11]<=32'b10111111110000100100000101101001;
        G_UP[12]<=32'b10111111110001000010001010010101;
        G_UP[13]<=32'b10000000000000000000000000000001;
        G_UP[14]<=32'b10000000000000000000000000000001;
        G_UP[15]<=32'b10000000000000000000000000000001;
        
        G_DOWN[0]<=32'b10000000000000000000000000000001;
        G_DOWN[1]<=32'b10000000000000000000000000000001;
        G_DOWN[2]<=32'b10000000000000000000000000000001;
        G_DOWN[3]<=32'b10111111110001000010000001100001;
        G_DOWN[4]<=32'b10111111110000100100000011110001;
        G_DOWN[5]<=32'b10111111110000111100000111111001;
        G_DOWN[6]<=32'b10111111110001011010001101101101;
        G_DOWN[7]<=32'b10111111110011111111001111111101;
        G_DOWN[8]<=32'b10111111110011111111000101101001;
        G_DOWN[9]<=32'b10111111110010100101001000000101;
        G_DOWN[10]<=32'b10111111110000111100000100001001;
        G_DOWN[11]<=32'b10000000000000000000000000000001;
        G_DOWN[12]<=32'b10000000000000000000000000000001;
        G_DOWN[13]<=32'b10000000000000000000000000000001;
        G_DOWN[14]<=32'b10000000000000000000000000000001;
        G_DOWN[15]<=32'b11111111111111111111111111111111;
            
        R_UP[0]<=32'b00000000000000000000000000000000;
        R_UP[1]<=32'b00000000000000000000000000000000;
        R_UP[2]<=32'b00000000000000000000000000000000;
        R_UP[3]<=32'b00000000000000000000000000000000;
        R_UP[4]<=32'b00000000000000000000000000000000;
        R_UP[5]<=32'b00000000000000000000000000000000;
        R_UP[6]<=32'b00000000000000000000000000000000;
        R_UP[7]<=32'b00000000000000000000000000000000;
        R_UP[8]<=32'b00000000000000000000000000000000;
        R_UP[9]<=32'b00000000000000000000000000000000;
        R_UP[10]<=32'b00000000000000000000000000000000;
        R_UP[11]<=32'b00000000000000000000000000000000;
        R_UP[12]<=32'b00000000000000000000000000000000;
        R_UP[13]<=32'b00000000000000000000000000000000;
        R_UP[14]<=32'b00000000000000000000000000000000;
        R_UP[15]<=32'b00000000000000000000000000000000;
        
        R_DOWN[0]<=32'b00000000000000000000000000000000;
        R_DOWN[1]<=32'b00000000000000000000000000000000;
        R_DOWN[2]<=32'b00000000000000000000000000000000;
        R_DOWN[3]<=32'b00000000000000000000000000000000;
        R_DOWN[4]<=32'b00000000000000000000000000000000;
        R_DOWN[5]<=32'b00000000000000000000000000000000;
        R_DOWN[6]<=32'b00000000000000000000000000000000;
        R_DOWN[7]<=32'b00000000000000000000000000000000;
        R_DOWN[8]<=32'b00000000000000000000000000000000;
        R_DOWN[9]<=32'b00000000000000000000000000000000;
        R_DOWN[10]<=32'b00000000000000000000000000000000;
        R_DOWN[11]<=32'b00000000000000000000000000000000;
        R_DOWN[12]<=32'b00000000000000000000000000000000;
        R_DOWN[13]<=32'b00000000000000000000000000000000;
        R_DOWN[14]<=32'b00000000000000000000000000000000;
        R_DOWN[15]<=32'b00000000000000000000000000000000;
            
		next_stage <= 3'b000;
		stage_select_flag <= 2'b0;
		count <= 0;
		
	end else if (cur_stage == OPENING ) begin //�I�[�v�j���O
	   
	   if(stage_select_flag == 2'b01) begin
	       if(sw3_raise == 1'b1)   next_stage <= 3'b001; 
	       else next_stage <= 3'b000;    
	   end else if(stage_select_flag == 2'b10) begin 
	       if(sw3_raise == 1'b1)   next_stage <= 3'b010; 
	       else next_stage <= 3'b000;     
	   end else if(stage_select_flag == 2'b11) begin
	       if(sw3_raise == 1'b1)   next_stage <= 3'b011; 
	       else next_stage <= 3'b000;  
	   end else    
	       next_stage <= 3'b000; 
      
	   if(sw2_raise == 1'b1) begin
	
	            stage_select_flag <= 2'b01;
                R_UP[0]<=32'b00000000000000000000000000000000;
                R_UP[1]<=32'b01111111111000000000000000000000;
                R_UP[2]<=32'b01111111111000000000000000000000;
                R_UP[3]<=32'b01111111111000000000000000000000;
                R_UP[4]<=32'b01111111111000000000000000000000;
                R_UP[5]<=32'b01111111111000000000000000000000;
                R_UP[6]<=32'b01111111111000000000000000000000;
                R_UP[7]<=32'b01111111111000000000000000000000;
                R_UP[8]<=32'b01111111111000000000000000000000;
                R_UP[9]<=32'b01111111111000000000000000000000;
                R_UP[10]<=32'b01111111111000000000000000000000;
                R_UP[11]<=32'b01111111111000000000000000000000;
                R_UP[12]<=32'b01111111111000000000000000000000;
                R_UP[13]<=32'b01111111111000000000000000000000;
                R_UP[14]<=32'b01111111111000000000000000000000;
                R_UP[15]<=32'b01111111111000000000000000000000;
                
                R_DOWN[0]<=32'b01111111111000000000000000000000;
                R_DOWN[1]<=32'b01111111111000000000000000000000;
                R_DOWN[2]<=32'b01111111111000000000000000000000;
                R_DOWN[3]<=32'b01111111111000000000000000000000;
                R_DOWN[4]<=32'b01111111111000000000000000000000;
                R_DOWN[5]<=32'b01111111111000000000000000000000;
                R_DOWN[6]<=32'b01111111111000000000000000000000;
                R_DOWN[7]<=32'b01111111111000000000000000000000;
                R_DOWN[8]<=32'b01111111111000000000000000000000;
                R_DOWN[9]<=32'b01111111111000000000000000000000;
                R_DOWN[10]<=32'b01111111111000000000000000000000;
                R_DOWN[11]<=32'b01111111111000000000000000000000;
                R_DOWN[12]<=32'b01111111111000000000000000000000;
                R_DOWN[13]<=32'b01111111111000000000000000000000;
                R_DOWN[14]<=32'b01111111111000000000000000000000;
                R_DOWN[15]<=32'b00000000000000000000000000000000;

    
	   end else if(sw1_raise == 1'b1) begin
	
	       stage_select_flag <= 2'b10;
            R_UP[0]<=32'b00000000000000000000000000000000;
            R_UP[1]<=32'b00000000000111111111100000000000;
            R_UP[2]<=32'b00000000000111111111100000000000;
            R_UP[3]<=32'b00000000000111111111100000000000;
            R_UP[4]<=32'b00000000000111111111100000000000;
            R_UP[5]<=32'b00000000000111111111100000000000;
            R_UP[6]<=32'b00000000000111111111100000000000;
            R_UP[7]<=32'b00000000000111111111100000000000;
            R_UP[8]<=32'b00000000000111111111100000000000;
            R_UP[9]<=32'b00000000000111111111100000000000;
            R_UP[10]<=32'b00000000000111111111100000000000;
            R_UP[11]<=32'b00000000000111111111100000000000;
            R_UP[12]<=32'b00000000000111111111100000000000;
            R_UP[13]<=32'b00000000000111111111100000000000;
            R_UP[14]<=32'b00000000000111111111100000000000;
            R_UP[15]<=32'b00000000000111111111100000000000;
            
            R_DOWN[0]<=32'b00000000000111111111100000000000;
            R_DOWN[1]<=32'b00000000000111111111100000000000;
            R_DOWN[2]<=32'b00000000000111111111100000000000;
            R_DOWN[3]<=32'b00000000000111111111100000000000;
            R_DOWN[4]<=32'b00000000000111111111100000000000;
            R_DOWN[5]<=32'b00000000000111111111100000000000;
            R_DOWN[6]<=32'b00000000000111111111100000000000;
            R_DOWN[7]<=32'b00000000000111111111100000000000;
            R_DOWN[8]<=32'b00000000000111111111100000000000;
            R_DOWN[9]<=32'b00000000000111111111100000000000;
            R_DOWN[10]<=32'b00000000000111111111100000000000;
            R_DOWN[11]<=32'b00000000000111111111100000000000;
            R_DOWN[12]<=32'b00000000000111111111100000000000;
            R_DOWN[13]<=32'b00000000000111111111100000000000;
            R_DOWN[14]<=32'b00000000000111111111100000000000;
            R_DOWN[15]<=32'b00000000000000000000000000000000;
    
	   end else if(sw0_raise == 1'b1) begin
	       stage_select_flag <= 2'b11;
            R_UP[0]<=32'b00000000000000000000000000000000;
            R_UP[1]<=32'b00000000000000000000011111111110;
            R_UP[2]<=32'b00000000000000000000011111111110;
            R_UP[3]<=32'b00000000000000000000011111111110;
            R_UP[4]<=32'b00000000000000000000011111111110;
            R_UP[5]<=32'b00000000000000000000011111111110;
            R_UP[6]<=32'b00000000000000000000011111111110;
            R_UP[7]<=32'b00000000000000000000011111111110;
            R_UP[8]<=32'b00000000000000000000011111111110;
            R_UP[9]<=32'b00000000000000000000011111111110;
            R_UP[10]<=32'b00000000000000000000011111111110;
            R_UP[11]<=32'b00000000000000000000011111111110;
            R_UP[12]<=32'b00000000000000000000011111111110;
            R_UP[13]<=32'b00000000000000000000011111111110;
            R_UP[14]<=32'b00000000000000000000011111111110;
            R_UP[15]<=32'b00000000000000000000011111111110;
            
            R_DOWN[0]<=32'b00000000000000000000011111111110;
            R_DOWN[1]<=32'b00000000000000000000011111111110;
            R_DOWN[2]<=32'b00000000000000000000011111111110;
            R_DOWN[3]<=32'b00000000000000000000011111111110;
            R_DOWN[4]<=32'b00000000000000000000011111111110;
            R_DOWN[5]<=32'b00000000000000000000011111111110;
            R_DOWN[6]<=32'b00000000000000000000011111111110;
            R_DOWN[7]<=32'b00000000000000000000011111111110;
            R_DOWN[8]<=32'b00000000000000000000011111111110;
            R_DOWN[9]<=32'b00000000000000000000011111111110;
            R_DOWN[10]<=32'b00000000000000000000011111111110;
            R_DOWN[11]<=32'b00000000000000000000011111111110;
            R_DOWN[12]<=32'b00000000000000000000011111111110;
            R_DOWN[13]<=32'b00000000000000000000011111111110;
            R_DOWN[14]<=32'b00000000000000000000011111111110;
            R_DOWN[15]<=32'b00000000000000000000000000000000;
       
	   end   
	   
	   
       if (count ==11999999) begin
            count <= 0;
            
            G_UP[0]<=32'b11111111111111111111111111111111;
            G_UP[1]<=32'b10000000000000000000000000000001;
            G_UP[2]<=32'b10000000000000000000000000000001;
            G_UP[3]<=32'b10000000000000000000000000000001;
            G_UP[4]<=32'b10000000000000000000000000000001;
            G_UP[5]<=32'b10111111110001000010000001100001;
            G_UP[6]<=32'b10111111110000100100000011110001;
            G_UP[7]<=32'b10111111110010111101000111111001;
            G_UP[8]<=32'b10111111110011011011001101101101;
            G_UP[9]<=32'b10111111110011111111001111111101;
            G_UP[10]<=32'b10111111110001111110000010010001;
            G_UP[11]<=32'b10111111110000100100000101101001;
            G_UP[12]<=32'b10111111110001000010001010010101;
            G_UP[13]<=32'b10000000000000000000000000000001;
            G_UP[14]<=32'b10000000000000000000000000000001;
            G_UP[15]<=32'b10000000000000000000000000000001;
            
            G_DOWN[0]<=32'b10000000000000000000000000000001;
            G_DOWN[1]<=32'b10000000000000000000000000000001;
            G_DOWN[2]<=32'b10000000000000000000000000000001;
            G_DOWN[3]<=32'b10111111110001000010000001100001;
            G_DOWN[4]<=32'b10111111110000100100000011110001;
            G_DOWN[5]<=32'b10111111110000111100000111111001;
            G_DOWN[6]<=32'b10111111110001011010001101101101;
            G_DOWN[7]<=32'b10111111110011111111001111111101;
            G_DOWN[8]<=32'b10111111110011111111000101101001;
            G_DOWN[9]<=32'b10111111110010100101001000000101;
            G_DOWN[10]<=32'b10111111110000111100000100001001;
            G_DOWN[11]<=32'b10000000000000000000000000000001;
            G_DOWN[12]<=32'b10000000000000000000000000000001;
            G_DOWN[13]<=32'b10000000000000000000000000000001;
            G_DOWN[14]<=32'b10000000000000000000000000000001;
            G_DOWN[15]<=32'b11111111111111111111111111111111;
    
    

        end else if (count==5999999) begin
        
        count <= count + 1;
        G_UP[0]<=32'b11111111111111111111111111111111;
        G_UP[1]<=32'b10000000000000000000000000000001;
        G_UP[2]<=32'b10000000000000000000000000000001;
        G_UP[3]<=32'b10000000000000000000000000000001;
        G_UP[4]<=32'b10000000000000000000000000000001;
        G_UP[5]<=32'b10111111110001000010000001100001;
        G_UP[6]<=32'b10111111110000100100000011110001;
        G_UP[7]<=32'b10111111110000111100000111111001;
        G_UP[8]<=32'b10111111110001011010001101101101;
        G_UP[9]<=32'b10111111110011111111001111111101;
        G_UP[10]<=32'b10111111110011111111000101101001;
        G_UP[11]<=32'b10111111110010100101001000000101;
        G_UP[12]<=32'b10111111110000111100000100001001;
        G_UP[13]<=32'b10000000000000000000000000000001;
        G_UP[14]<=32'b10000000000000000000000000000001;
        G_UP[15]<=32'b10000000000000000000000000000001;
        
        G_DOWN[0]<=32'b10000000000000000000000000000001;
        G_DOWN[1]<=32'b10000000000000000000000000000001;
        G_DOWN[2]<=32'b10000000000000000000000000000001;
        G_DOWN[3]<=32'b10111111110001000010000001100001;
        G_DOWN[4]<=32'b10111111110000100100000011110001;
        G_DOWN[5]<=32'b10111111110010111101000111111001;
        G_DOWN[6]<=32'b10111111110011011011001101101101;
        G_DOWN[7]<=32'b10111111110011111111001111111101;
        G_DOWN[8]<=32'b10111111110001111110000010010001;
        G_DOWN[9]<=32'b10111111110000100100000101101001;
        G_DOWN[10]<=32'b10111111110001000010001010010101;
        G_DOWN[11]<=32'b10000000000000000000000000000001;
        G_DOWN[12]<=32'b10000000000000000000000000000001;
        G_DOWN[13]<=32'b10000000000000000000000000000001;
        G_DOWN[14]<=32'b10000000000000000000000000000001;
        G_DOWN[15]<=32'b11111111111111111111111111111111;
        
    
    
        end else begin
          count <= count + 1;
          
       
       end
    end else if(cur_stage != OPENING ) begin //�I�[�v�j���O�X�e�[�W�łȂ���Ώ�����
        stage_select_flag <= 2'b00;
        R_UP[0]<=32'b00000000000000000000000000000000;
        R_UP[1]<=32'b00000000000000000000000000000000;
        R_UP[2]<=32'b00000000000000000000000000000000;
        R_UP[3]<=32'b00000000000000000000000000000000;
        R_UP[4]<=32'b00000000000000000000000000000000;
        R_UP[5]<=32'b00000000000000000000000000000000;
        R_UP[6]<=32'b00000000000000000000000000000000;
        R_UP[7]<=32'b00000000000000000000000000000000;
        R_UP[8]<=32'b00000000000000000000000000000000;
        R_UP[9]<=32'b00000000000000000000000000000000;
        R_UP[10]<=32'b00000000000000000000000000000000;
        R_UP[11]<=32'b00000000000000000000000000000000;
        R_UP[12]<=32'b00000000000000000000000000000000;
        R_UP[13]<=32'b00000000000000000000000000000000;
        R_UP[14]<=32'b00000000000000000000000000000000;
        R_UP[15]<=32'b00000000000000000000000000000000;
        
        R_DOWN[0]<=32'b00000000000000000000000000000000;
        R_DOWN[1]<=32'b00000000000000000000000000000000;
        R_DOWN[2]<=32'b00000000000000000000000000000000;
        R_DOWN[3]<=32'b00000000000000000000000000000000;
        R_DOWN[4]<=32'b00000000000000000000000000000000;
        R_DOWN[5]<=32'b00000000000000000000000000000000;
        R_DOWN[6]<=32'b00000000000000000000000000000000;
        R_DOWN[7]<=32'b00000000000000000000000000000000;
        R_DOWN[8]<=32'b00000000000000000000000000000000;
        R_DOWN[9]<=32'b00000000000000000000000000000000;
        R_DOWN[10]<=32'b00000000000000000000000000000000;
        R_DOWN[11]<=32'b00000000000000000000000000000000;
        R_DOWN[12]<=32'b00000000000000000000000000000000;
        R_DOWN[13]<=32'b00000000000000000000000000000000;
        R_DOWN[14]<=32'b00000000000000000000000000000000;
        R_DOWN[15]<=32'b00000000000000000000000000000000;
    
        
    end 
end


//�u�U�[�̐���
always @(posedge clk or posedge reset)begin
    if(reset == 1'b1) 
        sound_en <= 1'b0;
    else if(sw0_raise == 1'b1 |sw1_raise == 1'b1|sw2_raise == 1'b1) begin 
            sound_en <= 1'b1;       
    end else if( sound_count == BOM_SOUND ) begin
            sound_en <= 1'b0;
    end 
end


//�u�U�[���̒����J�E���g
always @(posedge clk or posedge reset)begin
    if(reset==1'b1)begin
        sound_count <=0;
    end else if(sound_en==1'b1) begin
        if (sound_count == BOM_SOUND) begin
            sound_count <= 0;
        end else if( sound_count < BOM_SOUND) begin    
            sound_count <= sound_count + 17'b1;
        end 
    end
end



endmodule





